
`define     BAGU_NOP                    2'h0

`define     BAGU_RLT                    2'h1
`define     BAGU_IMM                    2'h2
`define     BAGU_REG                    2'h3
