
`define     LSWIDTH_BYTE            2'b00
`define     LSWIDTH_HALF_WORD       2'b01
`define     LSWIDTH_WORD            2'b10
`define     LSWIDTH_DOUBLE_WORD     2'b11
