
`define     MUL_NOP                 1'b0
`define     MUL_EN                  1'b1