
module execute_mul_idffs (
    input   wire            clk,
    input   wire            resetn,

    //
    input   wire            i_valid,

    input   wire [31:0]     i_src0_value,
    input   wire [31:0]     i_src1_value,

    input   wire [3:0]      i_dst_rob,

    input   wire [7:0]      i_fid,

    input   wire [0:0]      i_mul_cmd,

    //
    output  wire            o_valid,

    output  wire [31:0]     o_src0_value,
    output  wire [31:0]     o_src1_value,

    output  wire [3:0]      o_dst_rob,

    output  wire [7:0]      o_fid,

    output  wire [0:0]      o_mul_cmd
);

    //
    reg         valid_R;

    reg [31:0]  src0_value_R;
    reg [31:0]  src1_value_R;

    reg [3:0]   dst_rob_R;

    reg [7:0]   fid_R;

    reg [0:0]   mul_cmd_R;

    always @(posedge clk) begin

        if (~resetn) begin
            valid_R <= 'b0;
        end
        else begin
            valid_R <= i_valid;
        end

        src0_value_R    <= i_src0_value;
        src1_value_R    <= i_src1_value;

        dst_rob_R       <= i_dst_rob;

        fid_R           <= i_fid;

        mul_cmd_R       <= i_mul_cmd;
    end

    //
    assign o_valid      = valid_R;
    
    assign o_src0_value = src0_value_R;
    assign o_src1_value = src1_value_R;

    assign o_dst_rob    = dst_rob_R;
    
    assign o_fid        = fid_R;

    assign o_mul_cmd    = mul_cmd_R;

    //

endmodule
