
module axi_constant32 (
    
);

endmodule
